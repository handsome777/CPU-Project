module InstructionMemory(Address, data);
	input [31:0] Address;
	output reg [31:0] data;

	reg [31:0] ROM[31:0]; //指令存储器的大小为2^32

	always @(*)
		case (Address[9:2])//9:2啥意思
0: data <=32'h08000003;
1: data <=32'h08000039;
2: data <=32'h08000038;
3: data <=32'h00008020;
4: data <=32'h3c104000;
5: data <=32'h22100018;
6: data <=32'h00008820;
7: data <=32'h3c110000;
8: data <=32'h22310002;
9: data <=32'h00002020;
10: data <=32'h00002820;
11: data <=32'h2210fff0;
12: data <=32'hae000000;
13: data <=32'h2210fff8;
14: data <=32'h2008fc18;
15: data <=32'hae080000;
16: data <=32'h2008ffff;
17: data <=32'h22100004;
18: data <=32'hae080000;
19: data <=32'h20080003;
20: data <=32'h22100004;
21: data <=32'hae080000;
22: data <=32'h22100018;
23: data <=32'h00001020;
24: data <=32'h8e080000;
25: data <=32'h01114824;
26: data <=32'h1120fffd;
27: data <=32'h2210fffc;
28: data <=32'h8e040000;
29: data <=32'h20860000;
30: data <=32'h22100004;
31: data <=32'h8e080000;
32: data <=32'h01114824;
33: data <=32'h1120fffd;
34: data <=32'h2210fffc;
35: data <=32'h8e050000;
36: data <=32'h20a70000;
37: data <=32'h22100004;
38: data <=32'h0800002d;
39: data <=32'h00805020;
40: data <=32'h01456022;
41: data <=32'h19800001;
42: data <=32'h01455022;
43: data <=32'h00a02020;
44: data <=32'h01402820;
45: data <=32'h1485fff9;
46: data <=32'h00801020;
47: data <=32'h3c104000;
48: data <=32'h2210000c;
49: data <=32'hae020000;
50: data <=32'h3c104000;
51: data <=32'h22100018;
52: data <=32'hae020000;
53: data <=32'h00001820;
54: data <=32'h00001820;
55: data <=32'h08000035;
56: data <=32'h03600008;
57: data <=32'h200dfff9;
58: data <=32'h0000b820;
59: data <=32'h3c174000;
60: data <=32'h22f70008;
61: data <=32'h8eee0000;
62: data <=32'h01ae6824;
63: data <=32'haeed0000;
64: data <=32'h22f7000c;
65: data <=32'h8eed0000;
66: data <=32'h31b60f00;
67: data <=32'h200e0100;
68: data <=32'h12c00007;
69: data <=32'h11d6000e;
70: data <=32'h000e7040;
71: data <=32'h11d60013;
72: data <=32'h000e7040;
73: data <=32'h11d60019;
74: data <=32'h000e7040;
75: data <=32'h11d60000;
76: data <=32'h00007820;
77: data <=32'h30ef00f0;
78: data <=32'h000f7902;
79: data <=32'h0c00006a;
80: data <=32'h20180100;
81: data <=32'h01f87825;
82: data <=32'haeef0000;
83: data <=32'h080000a9;
84: data <=32'h00007820;
85: data <=32'h30ef000f;
86: data <=32'h0c00006a;
87: data <=32'h20180200;
88: data <=32'h01f87825;
89: data <=32'haeef0000;
90: data <=32'h080000a9;
91: data <=32'h00007820;
92: data <=32'h30cf00f0;
93: data <=32'h000f7902;
94: data <=32'h0c00006a;
95: data <=32'h20180400;
96: data <=32'h01f87825;
97: data <=32'haeef0000;
98: data <=32'h080000a9;
99: data <=32'h00007820;
100: data <=32'h30cf000f;
101: data <=32'h0c00006a;
102: data <=32'h20180800;
103: data <=32'h01f87825;
104: data <=32'haeef0000;
105: data <=32'h080000a9;
106: data <=32'h200d0000;
107: data <=32'h15ed0002;
108: data <=32'h200f0040;
109: data <=32'h03e00008;
110: data <=32'h21ad0001;
111: data <=32'h15ed0002;
112: data <=32'h200f0079;
113: data <=32'h03e00008;
114: data <=32'h21ad0001;
115: data <=32'h15ed0002;
116: data <=32'h200f0024;
117: data <=32'h03e00008;
118: data <=32'h21ad0001;
119: data <=32'h15ed0002;
120: data <=32'h200f0030;
121: data <=32'h03e00008;
122: data <=32'h21ad0001;
123: data <=32'h15ed0002;
124: data <=32'h200f0019;
125: data <=32'h03e00008;
126: data <=32'h21ad0001;
127: data <=32'h15ed0002;
128: data <=32'h200f0012;
129: data <=32'h03e00008;
130: data <=32'h21ad0001;
131: data <=32'h15ed0002;
132: data <=32'h200f0002;
133: data <=32'h03e00008;
134: data <=32'h21ad0001;
135: data <=32'h15ed0002;
136: data <=32'h200f0078;
137: data <=32'h03e00008;
138: data <=32'h21ad0001;
139: data <=32'h15ed0002;
140: data <=32'h200f0000;
141: data <=32'h03e00008;
142: data <=32'h21ad0001;
143: data <=32'h15ed0002;
144: data <=32'h200f0010;
145: data <=32'h03e00008;
146: data <=32'h21ad0001;
147: data <=32'h15ed0002;
148: data <=32'h200f0008;
149: data <=32'h03e00008;
150: data <=32'h21ad0001;
151: data <=32'h15ed0002;
152: data <=32'h200f0003;
153: data <=32'h03e00008;
154: data <=32'h21ad0001;
155: data <=32'h15ed0002;
156: data <=32'h200f0046;
157: data <=32'h03e00008;
158: data <=32'h21ad0001;
159: data <=32'h15ed0002;
160: data <=32'h200f0021;
161: data <=32'h03e00008;
162: data <=32'h21ad0001;
163: data <=32'h15ed0002;
164: data <=32'h200f0006;
165: data <=32'h03e00008;
166: data <=32'h21ad0001;
167: data <=32'h200f000e;
168: data <=32'h03e00008;
169: data <=32'h0000b820;
170: data <=32'h3c174000;
171: data <=32'h22f70008;
172: data <=32'h8eee0000;
173: data <=32'h3c0f0000;
174: data <=32'h21ef0002;
175: data <=32'h01ee7025;
176: data <=32'haeee0000;
177: data <=32'h03400008;
			
			default: data <= 32'h80000000;
		endcase
		
endmodule